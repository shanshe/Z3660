localparam Z3660_VERS = 16'h0103;
localparam SYNTHESIS_VERS = 8'hAC;
localparam GPIO_VERS  = {SYNTHESIS_VERS,8'h00,Z3660_VERS};




